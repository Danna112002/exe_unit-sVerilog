`ifdef ALU_DEFINES
`define ALU_DEFINES

`define OPER_BITS       2
`define ALU_ADD        `OPER_BITS'd0
`define ALU_COMP       `OPER_BITS'd1
`define ALU_SET        `OPER_BITS'd2
`define ALU_CONV       `OPER_BITS'd3

`endif 